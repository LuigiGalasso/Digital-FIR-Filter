package CONSTANTS is
   constant NB : integer := 14;
   constant NT : integer := 9;
   --subtype coeff is array (0 to NT - 1) of std_logic_vector(NB - 1 downto 0);

end CONSTANTS;
